
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package test_data_pkg is
constant data_ch0 : unsigned(639 downto 0) := "0000000001111010000000000111101000000000011110010000000001111000000000000111100000000000011110110000000001111010000000000111101000000000011110110000000001111010000000000111100100000000100001100000000010100011000000001011111100000000110001000000000010111010000000001011000000000000101001000000000010011001000000001001001100000000100011000000000010001010000000001000010100000000100001100000000010000001000000001000000000000000011111110000000001111101000000000111101100000000011110100000000001111010000000000111100100000000011110000000000001111011000000000111101100000000011111010000000001111011000000000111110000000000011110000000000001111010";
constant data_ch1 : unsigned(639 downto 0) := "0000000101100101000000010110010000000001011001010000000101100101000000010110010000000001011010000000000101101000000000010110100000000001011010000000000101101000000000010110100000000001011101100000000110101000000000100001011100000010100001010000001010011101000000101000010100000010010101100000001000100111000000011111111100000001110111100000000111000101000000011010111100000001101000000000000110010011000000011000101100000001100001010000000101111101000000010111100100000001011101000000000101110001000000010110110100000001011010100000000101101011000000010110101000000001011010010000000101101000000000010110101000000001011001110000000101101000";
constant data_ch2 : unsigned(639 downto 0) := "0000000010001110000000001000111100000000100011100000000010001011000000001000101000000000100011010000000010001100000000001000101100000000100011000000000010001011000000001000101000000000100101010000000010101101000000001011101100000000101100100000000010100100000000001001111000000000100110000000000010010100000000001001010000000000100100100000000010010100000000001001001000000000100101010000000010010010000000001001000100000000100100010000000010001111000000001000111000000000100011100000000010001101000000001000110000000000100010100000000010001100000000001000110000000000100011010000000010001100000000001000111000000000100011000000000010001110";

end package;
